// sumador

module sum4(output wire[3:0] S, output wire c_out, input wire[3:0] A, input wire[3:0] B, input wire c_in);


  wire c1, c2, c3;
  fa b3(c_out, S[3], );
  fa b2();
  fa b1();
  fa b0();


endmodule